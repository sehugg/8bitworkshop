
`ifndef FONT_CP437_H
`define FONT_CP437_H

// PC font (code page 437)

module font_cp437_8x8(addr, data);

  input [10:0] addr;
  output [7:0] data;

  assign data = bitarray[addr];

  localparam [7:0] bitarray[0:2047] = '{
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00, //0
8'h7e,8'h81,8'ha5,8'h81,8'hbd,8'h99,8'h81,8'h7e, //1
8'h7e,8'hff,8'hdb,8'hff,8'hc3,8'he7,8'hff,8'h7e, //2
8'h6c,8'hfe,8'hfe,8'hfe,8'h7c,8'h38,8'h10,8'h00, //3
8'h10,8'h38,8'h7c,8'hfe,8'h7c,8'h38,8'h10,8'h00, //4
8'h38,8'h7c,8'h38,8'hfe,8'hfe,8'hd6,8'h10,8'h38, //5
8'h10,8'h10,8'h38,8'h7c,8'hfe,8'h7c,8'h10,8'h38, //6
8'h00,8'h00,8'h18,8'h3c,8'h3c,8'h18,8'h00,8'h00, //7
8'hff,8'hff,8'he7,8'hc3,8'hc3,8'he7,8'hff,8'hff, //8
8'h00,8'h3c,8'h66,8'h42,8'h42,8'h66,8'h3c,8'h00, //9
8'hff,8'hc3,8'h99,8'hbd,8'hbd,8'h99,8'hc3,8'hff, //10
8'h0f,8'h07,8'h0f,8'h7d,8'hcc,8'hcc,8'hcc,8'h78, //11
8'h3c,8'h66,8'h66,8'h66,8'h3c,8'h18,8'h7e,8'h18, //12
8'h3f,8'h33,8'h3f,8'h30,8'h30,8'h70,8'hf0,8'he0, //13
8'h7f,8'h63,8'h7f,8'h63,8'h63,8'h67,8'he6,8'hc0, //14
8'h99,8'h5a,8'h3c,8'he7,8'he7,8'h3c,8'h5a,8'h99, //15
8'h80,8'he0,8'hf8,8'hfe,8'hf8,8'he0,8'h80,8'h00, //16
8'h02,8'h0e,8'h3e,8'hfe,8'h3e,8'h0e,8'h02,8'h00, //17
8'h18,8'h3c,8'h7e,8'h18,8'h18,8'h7e,8'h3c,8'h18, //18
8'h66,8'h66,8'h66,8'h66,8'h66,8'h00,8'h66,8'h00, //19
8'h7f,8'hdb,8'hdb,8'h7b,8'h1b,8'h1b,8'h1b,8'h00, //20
8'h7e,8'hc3,8'h78,8'hcc,8'hcc,8'h78,8'h8c,8'hf8, //21
8'h00,8'h00,8'h00,8'h00,8'h7e,8'h7e,8'h7e,8'h00, //22
8'h18,8'h3c,8'h7e,8'h18,8'h7e,8'h3c,8'h18,8'hff, //23
8'h18,8'h3c,8'h7e,8'h18,8'h18,8'h18,8'h18,8'h00, //24
8'h18,8'h18,8'h18,8'h18,8'h7e,8'h3c,8'h18,8'h00, //25
8'h00,8'h18,8'h0c,8'hfe,8'h0c,8'h18,8'h00,8'h00, //26
8'h00,8'h30,8'h60,8'hfe,8'h60,8'h30,8'h00,8'h00, //27
8'h00,8'h00,8'hc0,8'hc0,8'hc0,8'hfe,8'h00,8'h00, //28
8'h00,8'h24,8'h66,8'hff,8'h66,8'h24,8'h00,8'h00, //29
8'h00,8'h18,8'h3c,8'h7e,8'hff,8'hff,8'h00,8'h00, //30
8'h00,8'hff,8'hff,8'h7e,8'h3c,8'h18,8'h00,8'h00, //31
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00, //32
8'h30,8'h78,8'h78,8'h30,8'h30,8'h00,8'h30,8'h00, //33
8'h6c,8'h6c,8'h6c,8'h00,8'h00,8'h00,8'h00,8'h00, //34
8'h6c,8'h6c,8'hfe,8'h6c,8'hfe,8'h6c,8'h6c,8'h00, //35
8'h30,8'h7c,8'hc0,8'h78,8'h0c,8'hf8,8'h30,8'h00, //36
8'h00,8'hc6,8'hcc,8'h18,8'h30,8'h66,8'hc6,8'h00, //37
8'h38,8'h6c,8'h38,8'h76,8'hdc,8'hcc,8'h76,8'h00, //38
8'h60,8'h60,8'hc0,8'h00,8'h00,8'h00,8'h00,8'h00, //39
8'h18,8'h30,8'h60,8'h60,8'h60,8'h30,8'h18,8'h00, //40
8'h60,8'h30,8'h18,8'h18,8'h18,8'h30,8'h60,8'h00, //41
8'h00,8'h66,8'h3c,8'hff,8'h3c,8'h66,8'h00,8'h00, //42
8'h00,8'h30,8'h30,8'hfc,8'h30,8'h30,8'h00,8'h00, //43
8'h00,8'h00,8'h00,8'h00,8'h00,8'h70,8'h30,8'h60, //44
8'h00,8'h00,8'h00,8'hfc,8'h00,8'h00,8'h00,8'h00, //45
8'h00,8'h00,8'h00,8'h00,8'h00,8'h30,8'h30,8'h00, //46
8'h06,8'h0c,8'h18,8'h30,8'h60,8'hc0,8'h80,8'h00, //47
8'h78,8'hcc,8'hdc,8'hfc,8'hec,8'hcc,8'h78,8'h00, //48
8'h30,8'hf0,8'h30,8'h30,8'h30,8'h30,8'hfc,8'h00, //49
8'h78,8'hcc,8'h0c,8'h38,8'h60,8'hcc,8'hfc,8'h00, //50
8'h78,8'hcc,8'h0c,8'h38,8'h0c,8'hcc,8'h78,8'h00, //51
8'h1c,8'h3c,8'h6c,8'hcc,8'hfe,8'h0c,8'h0c,8'h00, //52
8'hfc,8'hc0,8'hf8,8'h0c,8'h0c,8'hcc,8'h78,8'h00, //53
8'h38,8'h60,8'hc0,8'hf8,8'hcc,8'hcc,8'h78,8'h00, //54
8'hfc,8'hcc,8'h0c,8'h18,8'h30,8'h60,8'h60,8'h00, //55
8'h78,8'hcc,8'hcc,8'h78,8'hcc,8'hcc,8'h78,8'h00, //56
8'h78,8'hcc,8'hcc,8'h7c,8'h0c,8'h18,8'h70,8'h00, //57
8'h00,8'h00,8'h30,8'h30,8'h00,8'h30,8'h30,8'h00, //58
8'h00,8'h00,8'h30,8'h30,8'h00,8'h70,8'h30,8'h60, //59
8'h18,8'h30,8'h60,8'hc0,8'h60,8'h30,8'h18,8'h00, //60
8'h00,8'h00,8'hfc,8'h00,8'hfc,8'h00,8'h00,8'h00, //61
8'h60,8'h30,8'h18,8'h0c,8'h18,8'h30,8'h60,8'h00, //62
8'h78,8'hcc,8'h0c,8'h18,8'h30,8'h00,8'h30,8'h00, //63
8'h7c,8'hc6,8'hde,8'hde,8'hde,8'hc0,8'h78,8'h00, //64
8'h30,8'h78,8'hcc,8'hcc,8'hfc,8'hcc,8'hcc,8'h00, //65
8'hfc,8'h66,8'h66,8'h7c,8'h66,8'h66,8'hfc,8'h00, //66
8'h3c,8'h66,8'hc0,8'hc0,8'hc0,8'h66,8'h3c,8'h00, //67
8'hfc,8'h6c,8'h66,8'h66,8'h66,8'h6c,8'hfc,8'h00, //68
8'hfe,8'h62,8'h68,8'h78,8'h68,8'h62,8'hfe,8'h00, //69
8'hfe,8'h62,8'h68,8'h78,8'h68,8'h60,8'hf0,8'h00, //70
8'h3c,8'h66,8'hc0,8'hc0,8'hce,8'h66,8'h3e,8'h00, //71
8'hcc,8'hcc,8'hcc,8'hfc,8'hcc,8'hcc,8'hcc,8'h00, //72
8'h78,8'h30,8'h30,8'h30,8'h30,8'h30,8'h78,8'h00, //73
8'h1e,8'h0c,8'h0c,8'h0c,8'hcc,8'hcc,8'h78,8'h00, //74
8'he6,8'h66,8'h6c,8'h78,8'h6c,8'h66,8'he6,8'h00, //75
8'hf0,8'h60,8'h60,8'h60,8'h62,8'h66,8'hfe,8'h00, //76
8'hc6,8'hee,8'hfe,8'hd6,8'hc6,8'hc6,8'hc6,8'h00, //77
8'hc6,8'he6,8'hf6,8'hde,8'hce,8'hc6,8'hc6,8'h00, //78
8'h38,8'h6c,8'hc6,8'hc6,8'hc6,8'h6c,8'h38,8'h00, //79
8'hfc,8'h66,8'h66,8'h7c,8'h60,8'h60,8'hf0,8'h00, //80
8'h78,8'hcc,8'hcc,8'hcc,8'hdc,8'h78,8'h1c,8'h00, //81
8'hfc,8'h66,8'h66,8'h7c,8'h78,8'h6c,8'he6,8'h00, //82
8'h78,8'hcc,8'he0,8'h38,8'h1c,8'hcc,8'h78,8'h00, //83
8'hfc,8'hb4,8'h30,8'h30,8'h30,8'h30,8'h78,8'h00, //84
8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hfc,8'h00, //85
8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'h78,8'h30,8'h00, //86
8'hc6,8'hc6,8'hc6,8'hd6,8'hfe,8'hee,8'hc6,8'h00, //87
8'hc6,8'hc6,8'h6c,8'h38,8'h6c,8'hc6,8'hc6,8'h00, //88
8'hcc,8'hcc,8'hcc,8'h78,8'h30,8'h30,8'h78,8'h00, //89
8'hfe,8'hcc,8'h98,8'h30,8'h62,8'hc6,8'hfe,8'h00, //90
8'h78,8'h60,8'h60,8'h60,8'h60,8'h60,8'h78,8'h00, //91
8'hc0,8'h60,8'h30,8'h18,8'h0c,8'h06,8'h02,8'h00, //92
8'h78,8'h18,8'h18,8'h18,8'h18,8'h18,8'h78,8'h00, //93
8'h10,8'h38,8'h6c,8'hc6,8'h00,8'h00,8'h00,8'h00, //94
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff, //95
8'h30,8'h30,8'h18,8'h00,8'h00,8'h00,8'h00,8'h00, //96
8'h00,8'h00,8'h78,8'h0c,8'h7c,8'hcc,8'h76,8'h00, //97
8'he0,8'h60,8'h7c,8'h66,8'h66,8'h66,8'hbc,8'h00, //98
8'h00,8'h00,8'h78,8'hcc,8'hc0,8'hcc,8'h78,8'h00, //99
8'h1c,8'h0c,8'h0c,8'h7c,8'hcc,8'hcc,8'h76,8'h00, //100
8'h00,8'h00,8'h78,8'hcc,8'hfc,8'hc0,8'h78,8'h00, //101
8'h38,8'h6c,8'h60,8'hf0,8'h60,8'h60,8'hf0,8'h00, //102
8'h00,8'h00,8'h76,8'hcc,8'hcc,8'h7c,8'h0c,8'hf8, //103
8'he0,8'h60,8'h6c,8'h76,8'h66,8'h66,8'he6,8'h00, //104
8'h30,8'h00,8'h70,8'h30,8'h30,8'h30,8'h78,8'h00, //105
8'h18,8'h00,8'h78,8'h18,8'h18,8'h18,8'hd8,8'h70, //106
8'he0,8'h60,8'h66,8'h6c,8'h78,8'h6c,8'he6,8'h00, //107
8'h70,8'h30,8'h30,8'h30,8'h30,8'h30,8'h78,8'h00, //108
8'h00,8'h00,8'hec,8'hfe,8'hd6,8'hc6,8'hc6,8'h00, //109
8'h00,8'h00,8'hf8,8'hcc,8'hcc,8'hcc,8'hcc,8'h00, //110
8'h00,8'h00,8'h78,8'hcc,8'hcc,8'hcc,8'h78,8'h00, //111
8'h00,8'h00,8'hdc,8'h66,8'h66,8'h7c,8'h60,8'hf0, //112
8'h00,8'h00,8'h76,8'hcc,8'hcc,8'h7c,8'h0c,8'h1e, //113
8'h00,8'h00,8'hd8,8'h6c,8'h6c,8'h60,8'hf0,8'h00, //114
8'h00,8'h00,8'h7c,8'hc0,8'h78,8'h0c,8'hf8,8'h00, //115
8'h10,8'h30,8'h7c,8'h30,8'h30,8'h34,8'h18,8'h00, //116
8'h00,8'h00,8'hcc,8'hcc,8'hcc,8'hcc,8'h76,8'h00, //117
8'h00,8'h00,8'hcc,8'hcc,8'hcc,8'h78,8'h30,8'h00, //118
8'h00,8'h00,8'hc6,8'hc6,8'hd6,8'hfe,8'h6c,8'h00, //119
8'h00,8'h00,8'hc6,8'h6c,8'h38,8'h6c,8'hc6,8'h00, //120
8'h00,8'h00,8'hcc,8'hcc,8'hcc,8'h7c,8'h0c,8'hf8, //121
8'h00,8'h00,8'hfc,8'h98,8'h30,8'h64,8'hfc,8'h00, //122
8'h1c,8'h30,8'h30,8'he0,8'h30,8'h30,8'h1c,8'h00, //123
8'h18,8'h18,8'h18,8'h00,8'h18,8'h18,8'h18,8'h00, //124
8'he0,8'h30,8'h30,8'h1c,8'h30,8'h30,8'he0,8'h00, //125
8'h76,8'hdc,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00, //126
8'h10,8'h38,8'h6c,8'hc6,8'hc6,8'hc6,8'hfe,8'h00, //127
8'h78,8'hcc,8'hc0,8'hcc,8'h78,8'h18,8'h0c,8'h78, //128
8'h00,8'hcc,8'h00,8'hcc,8'hcc,8'hcc,8'h7e,8'h00, //129
8'h1c,8'h00,8'h78,8'hcc,8'hfc,8'hc0,8'h78,8'h00, //130
8'h7e,8'hc3,8'h3c,8'h06,8'h3e,8'h66,8'h3f,8'h00, //131
8'hcc,8'h00,8'h78,8'h0c,8'h7c,8'hcc,8'h7e,8'h00, //132
8'he0,8'h00,8'h78,8'h0c,8'h7c,8'hcc,8'h7e,8'h00, //133
8'h30,8'h30,8'h78,8'h0c,8'h7c,8'hcc,8'h7e,8'h00, //134
8'h00,8'h00,8'h7c,8'hc0,8'hc0,8'h7c,8'h06,8'h3c, //135
8'h7e,8'hc3,8'h3c,8'h66,8'h7e,8'h60,8'h3c,8'h00, //136
8'hcc,8'h00,8'h78,8'hcc,8'hfc,8'hc0,8'h78,8'h00, //137
8'he0,8'h00,8'h78,8'hcc,8'hfc,8'hc0,8'h78,8'h00, //138
8'hcc,8'h00,8'h70,8'h30,8'h30,8'h30,8'h78,8'h00, //139
8'h7c,8'hc6,8'h38,8'h18,8'h18,8'h18,8'h3c,8'h00, //140
8'he0,8'h00,8'h70,8'h30,8'h30,8'h30,8'h78,8'h00, //141
8'hcc,8'h30,8'h78,8'hcc,8'hcc,8'hfc,8'hcc,8'h00, //142
8'h30,8'h30,8'h00,8'h78,8'hcc,8'hfc,8'hcc,8'h00, //143
8'h1c,8'h00,8'hfc,8'h60,8'h78,8'h60,8'hfc,8'h00, //144
8'h00,8'h00,8'h7f,8'h0c,8'h7f,8'hcc,8'h7f,8'h00, //145
8'h3e,8'h6c,8'hcc,8'hfe,8'hcc,8'hcc,8'hce,8'h00, //146
8'h78,8'hcc,8'h00,8'h78,8'hcc,8'hcc,8'h78,8'h00, //147
8'h00,8'hcc,8'h00,8'h78,8'hcc,8'hcc,8'h78,8'h00, //148
8'h00,8'he0,8'h00,8'h78,8'hcc,8'hcc,8'h78,8'h00, //149
8'h78,8'hcc,8'h00,8'hcc,8'hcc,8'hcc,8'h7e,8'h00, //150
8'h00,8'he0,8'h00,8'hcc,8'hcc,8'hcc,8'h7e,8'h00, //151
8'h00,8'hcc,8'h00,8'hcc,8'hcc,8'hfc,8'h0c,8'hf8, //152
8'hc6,8'h38,8'h7c,8'hc6,8'hc6,8'h7c,8'h38,8'h00, //153
8'hcc,8'h00,8'hcc,8'hcc,8'hcc,8'hcc,8'h78,8'h00, //154
8'h18,8'h18,8'h7e,8'hc0,8'hc0,8'h7e,8'h18,8'h18, //155
8'h38,8'h6c,8'h64,8'hf0,8'h60,8'he6,8'hfc,8'h00, //156
8'hcc,8'hcc,8'h78,8'hfc,8'h30,8'hfc,8'h30,8'h00, //157
8'hf0,8'hd8,8'hd8,8'hf4,8'hcc,8'hde,8'hcc,8'h0e, //158
8'h0e,8'h1b,8'h18,8'h7e,8'h18,8'h18,8'hd8,8'h70, //159
8'h1c,8'h00,8'h78,8'h0c,8'h7c,8'hcc,8'h7e,8'h00, //160
8'h38,8'h00,8'h70,8'h30,8'h30,8'h30,8'h78,8'h00, //161
8'h00,8'h1c,8'h00,8'h78,8'hcc,8'hcc,8'h78,8'h00, //162
8'h00,8'h1c,8'h00,8'hcc,8'hcc,8'hcc,8'h7e,8'h00, //163
8'h00,8'hf8,8'h00,8'hf8,8'hcc,8'hcc,8'hcc,8'h00, //164
8'hfc,8'h00,8'hcc,8'hec,8'hfc,8'hdc,8'hcc,8'h00, //165
8'h3c,8'h6c,8'h6c,8'h3e,8'h00,8'h7e,8'h00,8'h00, //166
8'h3c,8'h66,8'h66,8'h3c,8'h00,8'h7e,8'h00,8'h00, //167
8'h30,8'h00,8'h30,8'h60,8'hc0,8'hcc,8'h78,8'h00, //168
8'h00,8'h00,8'h00,8'hfc,8'hc0,8'hc0,8'h00,8'h00, //169
8'h00,8'h00,8'h00,8'hfc,8'h0c,8'h0c,8'h00,8'h00, //170
8'hc6,8'hcc,8'hd8,8'h3e,8'h63,8'hce,8'h98,8'h1f, //171
8'hc6,8'hcc,8'hd8,8'hf3,8'h67,8'hcf,8'h9f,8'h03, //172
8'h00,8'h18,8'h00,8'h18,8'h18,8'h3c,8'h3c,8'h18, //173
8'h00,8'h33,8'h66,8'hcc,8'h66,8'h33,8'h00,8'h00, //174
8'h00,8'hcc,8'h66,8'h33,8'h66,8'hcc,8'h00,8'h00, //175
8'h22,8'h88,8'h22,8'h88,8'h22,8'h88,8'h22,8'h88, //176
8'h55,8'haa,8'h55,8'haa,8'h55,8'haa,8'h55,8'haa, //177
8'hdd,8'h77,8'hdd,8'h77,8'hdd,8'h77,8'hdd,8'h77, //178
8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18, //179
8'h18,8'h18,8'h18,8'h18,8'hf8,8'h18,8'h18,8'h18, //180
8'h18,8'h18,8'hf8,8'h18,8'hf8,8'h18,8'h18,8'h18, //181
8'h36,8'h36,8'h36,8'h36,8'hf6,8'h36,8'h36,8'h36, //182
8'h00,8'h00,8'h00,8'h00,8'hfe,8'h36,8'h36,8'h36, //183
8'h00,8'h00,8'hf8,8'h18,8'hf8,8'h18,8'h18,8'h18, //184
8'h36,8'h36,8'hf6,8'h06,8'hf6,8'h36,8'h36,8'h36, //185
8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36, //186
8'h00,8'h00,8'hfe,8'h06,8'hf6,8'h36,8'h36,8'h36, //187
8'h36,8'h36,8'hf6,8'h06,8'hfe,8'h00,8'h00,8'h00, //188
8'h36,8'h36,8'h36,8'h36,8'hfe,8'h00,8'h00,8'h00, //189
8'h18,8'h18,8'hf8,8'h18,8'hf8,8'h00,8'h00,8'h00, //190
8'h00,8'h00,8'h00,8'h00,8'hf8,8'h18,8'h18,8'h18, //191
8'h18,8'h18,8'h18,8'h18,8'h1f,8'h00,8'h00,8'h00, //192
8'h18,8'h18,8'h18,8'h18,8'hff,8'h00,8'h00,8'h00, //193
8'h00,8'h00,8'h00,8'h00,8'hff,8'h18,8'h18,8'h18, //194
8'h18,8'h18,8'h18,8'h18,8'h1f,8'h18,8'h18,8'h18, //195
8'h00,8'h00,8'h00,8'h00,8'hff,8'h00,8'h00,8'h00, //196
8'h18,8'h18,8'h18,8'h18,8'hff,8'h18,8'h18,8'h18, //197
8'h18,8'h18,8'h1f,8'h18,8'h1f,8'h18,8'h18,8'h18, //198
8'h36,8'h36,8'h36,8'h36,8'h37,8'h36,8'h36,8'h36, //199
8'h36,8'h36,8'h37,8'h30,8'h3f,8'h00,8'h00,8'h00, //200
8'h00,8'h00,8'h3f,8'h30,8'h37,8'h36,8'h36,8'h36, //201
8'h36,8'h36,8'hf7,8'h00,8'hff,8'h00,8'h00,8'h00, //202
8'h00,8'h00,8'hff,8'h00,8'hf7,8'h36,8'h36,8'h36, //203
8'h36,8'h36,8'h37,8'h30,8'h37,8'h36,8'h36,8'h36, //204
8'h00,8'h00,8'hff,8'h00,8'hff,8'h00,8'h00,8'h00, //205
8'h36,8'h36,8'hf7,8'h00,8'hf7,8'h36,8'h36,8'h36, //206
8'h18,8'h18,8'hff,8'h00,8'hff,8'h00,8'h00,8'h00, //207
8'h36,8'h36,8'h36,8'h36,8'hff,8'h00,8'h00,8'h00, //208
8'h00,8'h00,8'hff,8'h00,8'hff,8'h18,8'h18,8'h18, //209
8'h00,8'h00,8'h00,8'h00,8'hff,8'h36,8'h36,8'h36, //210
8'h36,8'h36,8'h36,8'h36,8'h3f,8'h00,8'h00,8'h00, //211
8'h18,8'h18,8'h1f,8'h18,8'h1f,8'h00,8'h00,8'h00, //212
8'h00,8'h00,8'h1f,8'h18,8'h1f,8'h18,8'h18,8'h18, //213
8'h00,8'h00,8'h00,8'h00,8'h3f,8'h36,8'h36,8'h36, //214
8'h36,8'h36,8'h36,8'h36,8'hf7,8'h36,8'h36,8'h36, //215
8'h18,8'h18,8'hff,8'h00,8'hff,8'h18,8'h18,8'h18, //216
8'h18,8'h18,8'h18,8'h18,8'hf8,8'h00,8'h00,8'h00, //217
8'h00,8'h00,8'h00,8'h00,8'h1f,8'h18,8'h18,8'h18, //218
8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff, //219
8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff, //220
8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0, //221
8'h0f,8'h0f,8'h0f,8'h0f,8'h0f,8'h0f,8'h0f,8'h0f, //222
8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00, //223
8'h00,8'h00,8'h76,8'hdc,8'hc8,8'hdc,8'h76,8'h00, //224
8'h00,8'h78,8'hcc,8'hf8,8'hcc,8'hf8,8'hc0,8'hc0, //225
8'h00,8'hfe,8'hc6,8'hc0,8'hc0,8'hc0,8'hc0,8'h00, //226
8'h00,8'hfe,8'h6c,8'h6c,8'h6c,8'h6c,8'h6c,8'h00, //227
8'hfe,8'h66,8'h30,8'h18,8'h30,8'h66,8'hfe,8'h00, //228
8'h00,8'h00,8'h7e,8'hcc,8'hcc,8'hcc,8'h78,8'h00, //229
8'h00,8'h66,8'h66,8'h66,8'h66,8'h7c,8'h60,8'hc0, //230
8'h00,8'h76,8'hdc,8'h18,8'h18,8'h18,8'h18,8'h00, //231
8'hfc,8'h30,8'h78,8'hcc,8'hcc,8'h78,8'h30,8'hfc, //232
8'h38,8'h6c,8'hc6,8'hfe,8'hc6,8'h6c,8'h38,8'h00, //233
8'h38,8'h6c,8'hc6,8'hc6,8'h6c,8'h6c,8'hee,8'h00, //234
8'h1c,8'h30,8'h18,8'h7c,8'hcc,8'hcc,8'h78,8'h00, //235
8'h00,8'h00,8'h7e,8'hdb,8'hdb,8'h7e,8'h00,8'h00, //236
8'h06,8'h0c,8'h7e,8'hdb,8'hdb,8'h7e,8'h60,8'hc0, //237
8'h3c,8'h60,8'hc0,8'hfc,8'hc0,8'h60,8'h3c,8'h00, //238
8'h78,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'h00, //239
8'h00,8'hfc,8'h00,8'hfc,8'h00,8'hfc,8'h00,8'h00, //240
8'h30,8'h30,8'hfc,8'h30,8'h30,8'h00,8'hfc,8'h00, //241
8'h60,8'h30,8'h18,8'h30,8'h60,8'h00,8'hfc,8'h00, //242
8'h18,8'h30,8'h60,8'h30,8'h18,8'h00,8'hfc,8'h00, //243
8'h0e,8'h1b,8'h1b,8'h18,8'h18,8'h18,8'h18,8'h18, //244
8'h18,8'h18,8'h18,8'h18,8'h18,8'hd8,8'hd8,8'h70, //245
8'h30,8'h30,8'h00,8'hfc,8'h00,8'h30,8'h30,8'h00, //246
8'h00,8'h72,8'h9c,8'h00,8'h72,8'h9c,8'h00,8'h00, //247
8'h38,8'h6c,8'h6c,8'h38,8'h00,8'h00,8'h00,8'h00, //248
8'h00,8'h00,8'h00,8'h18,8'h18,8'h00,8'h00,8'h00, //249
8'h00,8'h00,8'h00,8'h00,8'h18,8'h00,8'h00,8'h00, //250
8'h0f,8'h0c,8'h0c,8'h0c,8'hec,8'h6c,8'h3c,8'h1c, //251
8'h78,8'h6c,8'h6c,8'h6c,8'h6c,8'h00,8'h00,8'h00, //252
8'h78,8'h0c,8'h38,8'h60,8'h7c,8'h00,8'h00,8'h00, //253
8'h00,8'h00,8'h3c,8'h3c,8'h3c,8'h3c,8'h00,8'h00, //254
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00  //255
    };

endmodule

`endif
